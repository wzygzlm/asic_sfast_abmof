/usr/pack/global-28-kgf/dz/pdk/6U1x_2T8x_LB_2015.10/tech.lef