/usr/pack/global-28-kgf/arm/gf/cmos28slp/sc7mc_base_rvt_c34/r1p0/lef/sc7mc_cmos28slp_base_rvt_c34.lef