/usr/pack/global-28-kgf/arm/gf/cmos28lp/io_gppr_t18_mv11_mv18_tl25_rvt_dr/r6p0/lef/io_gppr_cmos28lp_t18_mv11_mv18_tl25_rvt_dr_6U1x_2T8x_LB.lef